-- ------------------------------------
library ieee ;
 use ieee . std_logic_1164 . all ;
 -- ------------------------------------
 entity Atividade2 is
 port (
 a , b , c, d: in bit ;
 s, t, u , v , w, x, y, z : out bit
 );
 end entity ;
 -- ------------------------------------
 architecture Atividade2 of Atividade2 is
 begin
	
 end architecture ;
-- ------------------------------------